`ifndef WDGRV_REGS_VH
`define WDGRV_REGS_VH
`define WDGRV_REGS_WDCSR_WDEN_BIT_WIDTH 1
`define WDGRV_REGS_WDCSR_WDEN_BIT_MASK 1'h1
`define WDGRV_REGS_WDCSR_WDEN_BIT_OFFSET 0
`define WDGRV_REGS_WDCSR_RVD1_BIT_WIDTH 1
`define WDGRV_REGS_WDCSR_RVD1_BIT_MASK 1'h1
`define WDGRV_REGS_WDCSR_RVD1_BIT_OFFSET 1
`define WDGRV_REGS_WDCSR_S1WTO_BIT_WIDTH 1
`define WDGRV_REGS_WDCSR_S1WTO_BIT_MASK 1'h1
`define WDGRV_REGS_WDCSR_S1WTO_BIT_OFFSET 2
`define WDGRV_REGS_WDCSR_S2WTO_BIT_WIDTH 1
`define WDGRV_REGS_WDCSR_S2WTO_BIT_MASK 1'h1
`define WDGRV_REGS_WDCSR_S2WTO_BIT_OFFSET 3
`define WDGRV_REGS_WDCSR_WTOCNT_BIT_WIDTH 10
`define WDGRV_REGS_WDCSR_WTOCNT_BIT_MASK 10'h3ff
`define WDGRV_REGS_WDCSR_WTOCNT_BIT_OFFSET 4
`define WDGRV_REGS_WDCSR_RVD2_BIT_WIDTH 18
`define WDGRV_REGS_WDCSR_RVD2_BIT_MASK 18'h3ffff
`define WDGRV_REGS_WDCSR_RVD2_BIT_OFFSET 14
`define WDGRV_REGS_WDCSR_BYTE_WIDTH 4
`define WDGRV_REGS_WDCSR_BYTE_SIZE 4
`define WDGRV_REGS_WDCSR_BYTE_OFFSET 3'h0
`define WDGRV_REGS_WDCNT_CNT_BIT_WIDTH 32
`define WDGRV_REGS_WDCNT_CNT_BIT_MASK 32'hffffffff
`define WDGRV_REGS_WDCNT_CNT_BIT_OFFSET 0
`define WDGRV_REGS_WDCNT_BYTE_WIDTH 4
`define WDGRV_REGS_WDCNT_BYTE_SIZE 4
`define WDGRV_REGS_WDCNT_BYTE_OFFSET 3'h4
`endif
