package wdgrv_regs_rtl_pkg;
  localparam int WDCSR_BYTE_WIDTH = 4;
  localparam int WDCSR_BYTE_SIZE = 4;
  localparam bit [2:0] WDCSR_BYTE_OFFSET = 3'h0;
  localparam int WDCSR_WDEN_BIT_WIDTH = 1;
  localparam bit WDCSR_WDEN_BIT_MASK = 1'h1;
  localparam int WDCSR_WDEN_BIT_OFFSET = 0;
  localparam int WDCSR_RVD1_BIT_WIDTH = 1;
  localparam bit WDCSR_RVD1_BIT_MASK = 1'h1;
  localparam int WDCSR_RVD1_BIT_OFFSET = 1;
  localparam int WDCSR_S1WTO_BIT_WIDTH = 1;
  localparam bit WDCSR_S1WTO_BIT_MASK = 1'h1;
  localparam int WDCSR_S1WTO_BIT_OFFSET = 2;
  localparam int WDCSR_S2WTO_BIT_WIDTH = 1;
  localparam bit WDCSR_S2WTO_BIT_MASK = 1'h1;
  localparam int WDCSR_S2WTO_BIT_OFFSET = 3;
  localparam int WDCSR_WTOCNT_BIT_WIDTH = 10;
  localparam bit [9:0] WDCSR_WTOCNT_BIT_MASK = 10'h3ff;
  localparam int WDCSR_WTOCNT_BIT_OFFSET = 4;
  localparam int WDCSR_RVD2_BIT_WIDTH = 18;
  localparam bit [17:0] WDCSR_RVD2_BIT_MASK = 18'h3ffff;
  localparam int WDCSR_RVD2_BIT_OFFSET = 14;
  localparam int WDCNT_BYTE_WIDTH = 4;
  localparam int WDCNT_BYTE_SIZE = 4;
  localparam bit [2:0] WDCNT_BYTE_OFFSET = 3'h4;
  localparam int WDCNT_CNT_BIT_WIDTH = 32;
  localparam bit [31:0] WDCNT_CNT_BIT_MASK = 32'hffffffff;
  localparam int WDCNT_CNT_BIT_OFFSET = 0;
endpackage
